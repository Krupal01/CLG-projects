*NMOS output characteristics
.model n1 NMOS(LEVEL=1 VTO=1V KP=20.179E-6 GAMMA=1.179
	+LAMBDA=0.005 PHI=0.66 uO=600 NSUB=5E15
	+Tox=1000E-8)
M_N 1 2 0 0 n1 w=2u l=2u
vgs 2 0 5v
vds 1 0 5v
.dc vds 0 5 0.1 vgs 0 5 1
.probe
.end

