// Copyright (C) 1991-2008 Altera Corporation
// Your use of Altera Corporation's design tools, logic functions 
// and other software and tools, and its AMPP partner logic 
// functions, and any output files from any of the foregoing 
// (including device programming or simulation files), and any 
// associated documentation or information are expressly subject 
// to the terms and conditions of the Altera Program License 
// Subscription Agreement, Altera MegaCore Function License 
// Agreement, or other applicable license agreement, including, 
// without limitation, that your use is for the sole purpose of 
// programming logic devices manufactured by Altera and sold by 
// Altera or its authorized distributors.  Please refer to the 
// applicable agreement for further details.

// PROGRAM		"Quartus II"
// VERSION		"Version 8.1 Build 163 10/28/2008 SJ Web Edition"
// CREATED ON	"Fri Oct 02 00:38:38 2020"

module Block1(
	pin_name,
	pin_name1,
	pin_name2,
	pin_name4
);


input	pin_name;
input	pin_name1;
input	pin_name2;
output	pin_name4;
reg	pin_name4;







endmodule
